library ieee;
use ieee.std_logic_1164.all;
Use ieee.numeric_std.all;
 
entity SR_FF is
	PORT( S,R,CLOCK: in std_logic;
			Q, QBAR: out std_logic);
end SR_FF;
 
Architecture behavioral of SR_FF is
begin
	PROCESS(CLOCK)
	variable tmp: std_logic;
	begin
	if(CLOCK='1' and CLOCK'EVENT) then
		if(S='0' and R='0')then
			tmp:=tmp;
		elsif(S='1' and R='1')then
			tmp:='Z';
		elsif(S='0' and R='1')then
			tmp:='0';
		else
			tmp:='1';
		end if;
	end if;
	Q <= tmp;
	QBAR <= not tmp;
	end PROCESS;
end behavioral;
